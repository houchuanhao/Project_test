library verilog;
use verilog.vl_types.all;
entity p1_vlg_tst is
end p1_vlg_tst;
